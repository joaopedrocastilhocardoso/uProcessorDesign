library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity StateMachine2Bits is
	port(
		clk, rst : in std_logic;
		state    : out unsigned(1 downto 0)
	);
	end entity;
	
architecture a_StateMachine2Bits of StateMachine2Bits is
	signal stateTemp : unsigned(1 downto 0) := "00";
	
	begin 
	
	process(clk, rst)
	begin
		if rst = '1' then -- if reset
			stateTemp <= "00";
			
		elsif rising_edge(clk) then 
			if stateTemp = "10" then -- if in stage 2 go back to stage 0
				stateTemp <= "00";
			else
				stateTemp <= 1 + stateTemp;
			end if;
		end if;
	end process;
	state <= stateTemp;
end architecture;